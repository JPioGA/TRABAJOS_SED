package tipos_esp is
generic ( MAX_ROUND : natrual := 99);
type natural_vector is array (0 to MAX_ROUND-1) of natural;

end tipos_esp;

package body tipos_esp is
end tipos_esp;