----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.12.2021 16:18:51
-- Design Name: 
-- Module Name: SIMON_DICE_TOP - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.tipos_esp.ALL;

entity SIMON_DICE_TOP is
--  Port ( );
end SIMON_DICE_TOP;

architecture structural of SIMON_DICE_TOP is

begin


end structural;
