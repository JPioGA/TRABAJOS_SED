----------------------------------------------------------------------------------
-- ENTIDAD TOP DEL JUEGO COMPLETO
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity DESCIFRA_EL_CODIGO_TOP is
    port (  CLK100MHZ   : in std_logic;
            CPU_RESETN  : in std_logic
    
    );
end DESCIFRA_EL_CODIGO_TOP;

architecture STRUCTURAL of DESCIFRA_EL_CODIGO_TOP is
    
begin


end STRUCTURAL;
