----------------------------------------------------------------------------------
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity USER_INPUT is
    Port ( CLK : in STD_LOGIC);
end USER_INPUT;

architecture Behavioral of USER_INPUT is

begin


end Behavioral;
