----------------------------------------------------------------------------------
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity FSM_1_SLAVE_INCHECK_TOP is
    port (
        CLK         : in std_logic;
        RST_N       : in std_logic
    );
end FSM_1_SLAVE_INCHECK_TOP;

architecture Behavioral of FSM_1_SLAVE_INCHECK_TOP is

begin


end Behavioral;
